library verilog;
use verilog.vl_types.all;
entity RTR_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end RTR_vlg_sample_tst;
