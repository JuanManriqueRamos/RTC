library verilog;
use verilog.vl_types.all;
entity RTR_vlg_vec_tst is
end RTR_vlg_vec_tst;
