library verilog;
use verilog.vl_types.all;
entity RTR is
    port(
        A0              : out    vl_logic;
        CLK             : in     vl_logic;
        B0              : out    vl_logic;
        C0              : out    vl_logic;
        D0              : out    vl_logic;
        E0              : out    vl_logic;
        F0              : out    vl_logic;
        G0              : out    vl_logic;
        B1              : out    vl_logic;
        C1              : out    vl_logic;
        D1              : out    vl_logic;
        E1              : out    vl_logic;
        F1              : out    vl_logic;
        G1              : out    vl_logic;
        A2              : out    vl_logic;
        B2              : out    vl_logic;
        C2              : out    vl_logic;
        D2              : out    vl_logic;
        F2              : out    vl_logic;
        G2              : out    vl_logic;
        A3              : out    vl_logic;
        B3              : out    vl_logic;
        C3              : out    vl_logic;
        D3              : out    vl_logic;
        E3              : out    vl_logic;
        F3              : out    vl_logic;
        G3              : out    vl_logic;
        A1              : out    vl_logic;
        E2              : out    vl_logic
    );
end RTR;
